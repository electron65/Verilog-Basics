`timescale 1ns/1n

module not_gate(a,x);

input a;
output x;

not U1(x, a);

endmodule
