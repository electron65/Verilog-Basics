`timescale 1ns/1ns

module not_prim(a,x);

input a;
output x;

not U1(x, a);

endmodule
