module notgate(input a,
		output x
		); // define the module, definition of input and output

assign x = ~a;

endmodule // end module
